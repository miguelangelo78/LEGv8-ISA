/****************************************************************************
 * pipeline_buffers.sv
 ****************************************************************************/

/**
 * Module: Pipes
 * 
 * TODO: Add module documentation
 */
module Pipes;

endmodule
