/****************************************************************************
 * legv8.sv
 ****************************************************************************/
`include "microcode.sv"

/**
 * Module: legv8
 * 
 * TODO: Add module documentation
 */
module LEGv8(input clk, input restart_cpu);
 	
endmodule